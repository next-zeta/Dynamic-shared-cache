module comparator_port (
    input  [4:0] port,
    input  [10:0] a,  
    input  [10:0] b,  
    input  [10:0] c,  
    output [4:0] port_max  
);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
// 中间信号用于存储比较结果
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
    logic [10:0] max_ab;
    logic [4:0]  max_tmp;
    logic [10:0] max_bc;
    logic [4:0]  max;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
// 比较a和b的大小
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        if (a > b) begin
            max_ab <= a;
            max_tmp <= port - 7;
        end
        else begin
            max_ab = b;
            max_tmp <= port;
        end
    end

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
// 比较max_ab和c的大小
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always_comb begin
        if (max_ab > c) begin
            max <= max_tmp;
        end
        else begin
            max <= port + 7;
        end
    end

    assign port_max = max;

endmodule
