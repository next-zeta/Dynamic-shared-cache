module bitmap(
    input logic clk,
    input logic rst_n,
    
);